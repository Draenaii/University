skyddet av miljön . Därför förespråkar vi att man fastslår en politik för jordbruket och landsbygdens utveckling som överensstämmer med de mål som vi har satt upp och att landsbygden
