effektivitet , som kan användas till vad som helst ,
