historiska arvet hade också skadats , vilket det sorgliga exemplet Versailles slottspark vittnar om . Inför en sådan katastrof förefaller det därför naturligt att den nationella och europeiska solidariteten kommer de olycksdrabbade och de mest berörda personerna till del . Men i likhet med vad föregående talare har sagt , och vad ni , herr kommissionär , svarade min kollega Jean-Claude Martinez angående en annan tragedi - nämligen översvämningarna i sydvästra Frankrike i november månad - är det visserligen så att ni ser med oro på katastroferna , men det
