stor vikt . På den punkten är förslaget helt enkelt
