mot naziregimen . ( Applåder ) Herr Poettering ! Jag ifrågasätter inte er demokratiska oro , men jag tror att ni begår ett allvarligt politiskt misstag . Och för att parafrasera en av mina ryktbara landsmän , Europas fader , Paul-Henri Spaak , skall jag säga att för er del är det inte för sent , men det är dags att ändra åsikt . Fru talman ! I dag ställs Europeiska unionen enligt min grupp inför sin största politiska och etiska utmaning sedan den bildades . Unionen har förvisso upplevt
