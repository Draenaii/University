, de mål , mekanismer och lagbestämmelser som berör sektorn , så stöder vi dem till fullo . Beslutar sig kommissionen för att driva igenom dessa informativa bemödanden så skulle inget , ärade kollegor , göra oss gladare . Vid kommissionärens sista inställelse inför kommissionen erkände han att det var absolut nödvändigt . Fischler sade att vi har problem med marketing och att det är nödvändigt att informera och värna om vår modell . Intern information - mot den egna sektorn , inom vilken man ofta inte känner till eller
