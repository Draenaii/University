måste ställas inför rätta . Att rädda och skydda liv under dessa extraordinära omständigheter utgör en oskiljaktig del av den humanitära rätten . ECHO : s roll i Colombia ,
