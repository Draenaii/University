. Jag frågar ju inte detta utan orsak . Ni har med all rätt sagt att försiktighetsprincipen är nödvändig just när vetenskapen ännu inte har några bevis . Hur skall
