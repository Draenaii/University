insatser . Hur som helst vill jag meddela parlamentet att en särskild delegation från kommissionen kommer att ge sig av för att granska sällskapet RINA den 28 : e nästa
