en rättvis territorialpolitik . I riktlinjerna tas hänsyn till två horisontella principer : landsbygdsutveckling och , fru föredragande , jag innefattar i landsbygdsutveckling också frågan om hållbara transporter som jag personligen fäster stor betydelse vid sedan länge - bl.a. när jag tänker på min tid som miljöminister i mitt land - och den andra principen handlar om lika möjligheter , framför allt för män och kvinnor , liksom den europeiska strategin för sysselsättning och ramen för den ekonomiska och monetära unionen . Avslutningsvis och för att bemöta den oro ni
