att vi anser , och det framgår av ordalydelsen i
