- i varje fall delvis - en ny kommission .
